magic
tech sky130A
magscale 1 2
timestamp 1713724750
<< error_s >>
rect 5151 -502 6458 -251
rect 5151 -1140 5384 -502
rect 6376 -1140 6458 -502
rect 5151 -2113 5437 -1140
rect 6172 -2113 6458 -1140
rect 5151 -2399 6458 -2113
<< dnwell >>
rect 5231 -2319 6378 -331
<< locali >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 2319 -509 3279 -340
rect 5238 -369 6341 -340
rect 5238 -492 5459 -369
rect 6304 -492 6341 -369
rect 5238 -538 6341 -492
rect 5238 -1104 5421 -538
rect 5237 -1740 5421 -1226
rect 1183 -2314 2143 -1781
rect 5554 -2034 6341 -1774
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5237 -2121 6341 -2034
rect 5237 -2244 5279 -2121
rect 6279 -2244 6341 -2121
rect 5237 -2314 6341 -2244
<< viali >>
rect 1223 -493 2106 -370
rect 5459 -492 6304 -369
rect 2357 -2286 3240 -2163
rect 5279 -2244 6279 -2121
<< metal1 >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 5421 -369 6341 -340
rect 5421 -492 5459 -369
rect 6304 -492 6341 -369
rect 5421 -538 6341 -492
rect 1183 -758 1325 -539
rect 1353 -710 1363 -658
rect 1963 -710 1973 -658
rect 2489 -670 2499 -618
rect 3099 -670 3109 -618
rect 1183 -959 1357 -758
rect 1969 -830 2494 -746
rect 1969 -887 2205 -830
rect 2345 -887 2494 -830
rect 1969 -958 2494 -887
rect 1183 -1362 1325 -959
rect 1353 -1058 1363 -1006
rect 1963 -1058 1973 -1006
rect 2489 -1167 2505 -1151
rect 3095 -1167 3105 -1151
rect 2489 -1219 2499 -1167
rect 3099 -1219 3105 -1167
rect 1353 -1314 1363 -1262
rect 1963 -1314 1973 -1262
rect 1183 -1562 1357 -1362
rect 1969 -1427 2461 -1362
rect 1969 -1484 1985 -1427
rect 2125 -1484 2461 -1427
rect 2489 -1457 2499 -1405
rect 3099 -1457 3105 -1405
rect 2489 -1473 2504 -1457
rect 3095 -1473 3105 -1457
rect 1969 -1562 2461 -1484
rect 2462 -1562 2493 -1505
rect 1353 -1662 1363 -1610
rect 1963 -1662 1973 -1610
rect 2271 -1905 2493 -1562
rect 2489 -1953 3109 -1937
rect 2489 -2005 2499 -1953
rect 3099 -2005 3109 -1953
rect 3137 -2115 3279 -718
rect 5421 -721 5543 -538
rect 5571 -673 5581 -621
rect 6181 -673 6191 -621
rect 5421 -921 5575 -721
rect 6187 -921 6341 -721
rect 5571 -1021 5581 -969
rect 6181 -1021 6188 -969
rect 6216 -1104 6341 -921
rect 5455 -1225 6341 -1104
rect 5455 -1226 6307 -1225
rect 5455 -1400 5546 -1226
rect 5574 -1352 5580 -1300
rect 6181 -1352 6191 -1300
rect 5574 -1368 6191 -1352
rect 5455 -1599 5523 -1400
rect 5575 -1599 5585 -1400
rect 5455 -1600 5574 -1599
rect 6187 -1600 6341 -1400
rect 5571 -1700 5581 -1648
rect 6182 -1700 6192 -1648
rect 5330 -1926 5339 -1848
rect 5479 -1926 5489 -1848
rect 6220 -2034 6341 -1600
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5237 -2121 6341 -2034
rect 5237 -2244 5279 -2121
rect 6279 -2244 6341 -2121
rect 5237 -2314 6341 -2244
<< via1 >>
rect 1363 -710 1963 -658
rect 2499 -670 3099 -618
rect 2205 -887 2345 -830
rect 1363 -1058 1963 -1006
rect 2499 -1219 3099 -1167
rect 1363 -1314 1963 -1262
rect 1985 -1484 2125 -1427
rect 2499 -1457 3099 -1405
rect 1363 -1662 1963 -1610
rect 2499 -2005 3099 -1953
rect 5581 -673 6181 -621
rect 5581 -1021 6181 -969
rect 5580 -1352 6181 -1300
rect 5523 -1599 5575 -1400
rect 5581 -1700 6182 -1648
rect 5339 -1926 5479 -1848
<< metal2 >>
rect 2499 -616 6181 -606
rect 2499 -618 5342 -616
rect 1363 -657 2135 -643
rect 1363 -658 1985 -657
rect 1963 -710 1985 -658
rect 1363 -714 1985 -710
rect 2125 -714 2135 -657
rect 3099 -670 5342 -618
rect 2499 -673 5342 -670
rect 5482 -621 6181 -616
rect 5482 -673 5581 -621
rect 2499 -683 6181 -673
rect 1363 -720 2135 -714
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -897 2355 -887
rect 5330 -969 6181 -959
rect 1363 -1006 2135 -996
rect 1963 -1058 1985 -1006
rect 1363 -1063 1985 -1058
rect 2125 -1063 2135 -1006
rect 5330 -1026 5340 -969
rect 5480 -1021 5581 -969
rect 5480 -1026 6181 -1021
rect 5330 -1036 6181 -1026
rect 1363 -1068 2135 -1063
rect 1363 -1073 2125 -1068
rect 2499 -1164 5490 -1157
rect 2499 -1167 5340 -1164
rect 3099 -1219 5340 -1167
rect 2499 -1221 5340 -1219
rect 5480 -1221 5490 -1164
rect 2499 -1229 5490 -1221
rect 1363 -1257 2355 -1247
rect 1363 -1262 2205 -1257
rect 1963 -1314 2205 -1262
rect 2345 -1314 2355 -1257
rect 1363 -1324 2355 -1314
rect 5330 -1294 6181 -1285
rect 5330 -1351 5340 -1294
rect 5480 -1300 6181 -1294
rect 5480 -1351 5580 -1300
rect 5330 -1352 5580 -1351
rect 5330 -1362 6181 -1352
rect 2499 -1400 5575 -1390
rect 2499 -1405 3177 -1400
rect 1975 -1427 2135 -1417
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 3099 -1457 3177 -1405
rect 3317 -1457 5523 -1400
rect 2499 -1467 5523 -1457
rect 1975 -1494 2135 -1484
rect 1363 -1610 2355 -1600
rect 5523 -1609 5575 -1599
rect 1963 -1662 2205 -1610
rect 1363 -1667 2205 -1662
rect 2345 -1667 2355 -1610
rect 1363 -1672 2355 -1667
rect 5330 -1648 6182 -1638
rect 5330 -1705 5340 -1648
rect 5480 -1700 5581 -1648
rect 5480 -1705 6182 -1700
rect 5330 -1715 6182 -1705
rect 5339 -1848 5479 -1838
rect 5339 -1936 5479 -1926
rect 2499 -1952 3327 -1943
rect 2499 -1953 3177 -1952
rect 3099 -2005 3177 -1953
rect 2499 -2009 3177 -2005
rect 3317 -2009 3327 -1952
rect 2499 -2015 3327 -2009
<< via2 >>
rect 1985 -714 2125 -657
rect 5342 -673 5482 -616
rect 2205 -887 2345 -830
rect 1985 -1063 2125 -1006
rect 5340 -1026 5480 -969
rect 5340 -1221 5480 -1164
rect 2205 -1314 2345 -1257
rect 5340 -1351 5480 -1294
rect 1985 -1484 2125 -1427
rect 3177 -1457 3317 -1400
rect 2205 -1667 2345 -1610
rect 5340 -1705 5480 -1648
rect 5339 -1926 5479 -1848
rect 3177 -2009 3317 -1952
<< metal3 >>
rect 5330 -616 5491 -606
rect 1975 -657 2135 -648
rect 1975 -714 1985 -657
rect 2125 -714 2135 -657
rect 1975 -1006 2135 -714
rect 5330 -673 5342 -616
rect 5482 -673 5491 -616
rect 1975 -1063 1985 -1006
rect 2125 -1063 2135 -1006
rect 1975 -1427 2135 -1063
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 1975 -1494 2135 -1484
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -1257 2355 -887
rect 2195 -1314 2205 -1257
rect 2345 -1314 2355 -1257
rect 2195 -1610 2355 -1314
rect 5330 -969 5491 -673
rect 5330 -1026 5340 -969
rect 5480 -1026 5491 -969
rect 5330 -1164 5491 -1026
rect 5330 -1221 5340 -1164
rect 5480 -1221 5491 -1164
rect 5330 -1294 5491 -1221
rect 5330 -1351 5340 -1294
rect 5480 -1351 5491 -1294
rect 2195 -1667 2205 -1610
rect 2345 -1667 2355 -1610
rect 2195 -1672 2355 -1667
rect 3167 -1400 3327 -1390
rect 3167 -1457 3177 -1400
rect 3317 -1457 3327 -1400
rect 3167 -1952 3327 -1457
rect 3167 -2009 3177 -1952
rect 3317 -2009 3327 -1952
rect 3167 -2014 3327 -2009
rect 5330 -1648 5491 -1351
rect 5330 -1705 5340 -1648
rect 5480 -1705 5491 -1648
rect 5330 -1848 5491 -1705
rect 5330 -1926 5339 -1848
rect 5479 -1926 5491 -1848
rect 5330 -2015 5491 -1926
use sky130_fd_pr__diode_pw2nd_05v5_37RBXE  sky130_fd_pr__diode_pw2nd_05v5_37RBXE_0 paramcells
timestamp 1713221383
transform 0 1 5408 -1 0 -1887
box -183 -208 183 208
use sky130_fd_pr__nfet_01v8_MG6U6H  sky130_fd_pr__nfet_01v8_MG6U6H_0 paramcells
timestamp 1713221383
transform 1 0 5880 0 1 -1500
box -496 -310 496 310
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0 paramcells
timestamp 1713228232
transform -1 0 2799 0 1 -1705
box -528 -458 528 458
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1
timestamp 1713228232
transform -1 0 2799 0 1 -919
box -528 -458 528 458
use sky130_fd_pr__pfet_01v8_J2L9Q3  sky130_fd_pr__pfet_01v8_J2L9Q3_0 paramcells
timestamp 1713221383
transform 1 0 5880 0 1 -821
box -496 -319 496 319
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0 paramcells
timestamp 1713221383
transform 1 0 1663 0 -1 -1462
box -558 -397 558 397
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1
timestamp 1713221383
transform 1 0 1663 0 -1 -858
box -558 -397 558 397
<< labels >>
flabel space 1105 -1255 2221 -461 0 FreeSans 1600 0 0 0 M3
flabel space 2271 -1377 3327 -461 0 FreeSans 1600 0 0 0 M5
flabel space 2271 -2163 3327 -1247 0 FreeSans 1600 0 0 0 M6
flabel metal1 1183 -539 2143 -340 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 1363 -1662 1963 -1610 0 FreeSans 800 0 0 0 out_b
port 5 nsew
flabel metal2 1363 -710 1963 -658 0 FreeSans 800 0 0 0 out
port 4 nsew
flabel space 1105 -1859 2221 -1065 0 FreeSans 1600 0 0 0 M4
flabel metal2 3317 -1467 3773 -1390 0 FreeSans 800 0 0 0 in_b
flabel metal1 2319 -2314 3279 -2115 0 FreeSans 1600 0 0 0 avss
port 6 nsew
flabel metal3 5330 -2015 5491 -1926 0 FreeSans 1600 0 0 0 in
port 3 nsew
flabel metal1 5237 -2313 6341 -2244 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
flabel space 5384 -1140 6376 -502 0 FreeSans 1600 0 0 0 M2
flabel space 5384 -1810 6376 -1190 0 FreeSans 1600 0 0 0 M1
flabel metal1 5421 -409 6341 -340 0 FreeSans 1600 0 0 0 dvdd
port 2 nsew
<< end >>
