magic
tech sky130A
magscale 1 2
timestamp 1726593208
<< pwell >>
rect -1259 717 12781 18089
rect -1259 -369 12733 717
rect -1259 -399 13789 -369
<< mvpsubdiff >>
rect -1193 18011 12715 18023
rect -1193 17977 -1085 18011
rect 12607 17977 12715 18011
rect -1193 17965 12715 17977
rect -1193 17915 -1135 17965
rect -1193 -225 -1181 17915
rect -1147 -225 -1135 17915
rect -1193 -275 -1135 -225
rect 12657 17915 12715 17965
rect 12657 -225 12669 17915
rect 12703 -225 12715 17915
rect 12657 -275 12715 -225
rect -1193 -287 12715 -275
rect -1193 -321 -1085 -287
rect 12607 -321 12715 -287
rect -1193 -333 12715 -321
<< mvpsubdiffcont >>
rect -1085 17977 12607 18011
rect -1181 -225 -1147 17915
rect 12669 -225 12703 17915
rect -1085 -321 12607 -287
<< locali >>
rect -1259 18011 12781 18089
rect -1259 17977 -1085 18011
rect 12607 17977 12781 18011
rect -1259 17932 12781 17977
rect -1259 17915 -1102 17932
rect -1259 -225 -1181 17915
rect -1147 -225 -1102 17915
rect -1259 -242 -1102 -225
rect 12624 17915 12781 17932
rect 12624 -225 12669 17915
rect 12703 747 12781 17915
rect 12703 653 14153 747
rect 12703 -225 12827 653
rect 12624 -242 12827 -225
rect -1259 -275 12827 -242
rect 13695 327 14153 653
rect 13695 51 13857 327
rect 14083 51 14153 327
rect 13695 -67 14153 51
rect 13695 -275 13860 -67
rect -1259 -287 13860 -275
rect -1259 -321 -1085 -287
rect 12607 -321 13860 -287
rect -1259 -791 13860 -321
rect -1259 -1191 -357 -791
rect 14080 -1191 14153 -67
rect -1259 -1438 14153 -1191
<< viali >>
rect 13860 -791 14080 -67
rect -357 -1191 14080 -791
<< metal1 >>
rect -1259 19108 12781 19128
rect -1259 18253 10921 19108
rect 11333 18253 12781 19108
rect -1259 18233 12781 18253
rect -1039 17587 12561 17869
rect -1039 103 75 17587
rect 10911 17491 11343 17501
rect 179 16831 611 17491
rect 3399 17209 4367 17491
rect 7155 17209 8123 17491
rect 10911 17199 11343 17209
rect 179 16075 611 16735
rect 3399 16453 3831 17113
rect 3935 16453 4367 17113
rect 7155 16831 8123 17113
rect 179 15319 611 15979
rect 3399 15697 3831 16357
rect 3935 15697 4367 16357
rect 7155 16075 7587 16735
rect 7691 16075 8123 16735
rect 10911 16453 11343 17113
rect 179 14563 611 15223
rect 3399 14941 3831 15601
rect 3935 14941 4367 15601
rect 7155 15319 7587 15979
rect 7691 15319 8123 15979
rect 10911 15697 11343 16357
rect 179 13807 611 14467
rect 3399 14185 3831 14845
rect 3935 14185 4367 14845
rect 7155 14563 7587 15223
rect 7691 14563 8123 15223
rect 10911 14941 11343 15601
rect 179 13051 611 13711
rect 3399 13429 3831 14089
rect 3935 13429 4367 14089
rect 7155 13807 7587 14467
rect 7691 13807 8123 14467
rect 10911 14185 11343 14845
rect 179 12295 611 12955
rect 3399 12673 3831 13333
rect 3935 12673 4367 13333
rect 7155 13051 7587 13711
rect 7691 13051 8123 13711
rect 10911 13429 11343 14089
rect 179 11539 611 12199
rect 3399 11917 3831 12577
rect 3935 11917 4367 12577
rect 7155 12295 7587 12955
rect 7691 12295 8123 12955
rect 10911 12673 11343 13333
rect 179 10783 611 11443
rect 3399 11161 3831 11821
rect 3935 11161 4367 11821
rect 7155 11539 7587 12199
rect 7691 11539 8123 12199
rect 10911 11917 11343 12577
rect 10911 11443 11343 11821
rect 179 10027 611 10687
rect 3399 10405 3831 11065
rect 3935 10405 4367 11065
rect 7155 10783 7587 11443
rect 7691 10783 8123 11443
rect 10901 11161 10911 11443
rect 11343 11161 11353 11443
rect 10911 10687 11343 11065
rect 179 9271 611 9931
rect 3399 9649 3831 10309
rect 3935 9649 4367 10309
rect 7155 10027 7587 10687
rect 7691 10027 8123 10687
rect 10901 10405 10911 10687
rect 11343 10405 11353 10687
rect 10911 9931 11343 10309
rect 179 8515 611 9175
rect 3399 8893 3831 9553
rect 3935 8893 4367 9553
rect 7155 9271 7587 9931
rect 7691 9271 8123 9931
rect 10901 9649 10911 9931
rect 11343 9649 11353 9931
rect 10911 9175 11343 9553
rect 179 7759 611 8419
rect 3399 8137 3831 8797
rect 3935 8137 4367 8797
rect 7155 8515 7587 9175
rect 7691 8797 8123 9175
rect 10901 8893 10911 9175
rect 11343 8893 11353 9175
rect 7681 8515 7691 8797
rect 8123 8515 8133 8797
rect 10911 8419 11343 8797
rect 179 7003 611 7663
rect 3399 7381 3831 8041
rect 3935 7381 4367 8041
rect 7155 7759 7587 8419
rect 7691 8041 8123 8419
rect 10901 8137 11353 8419
rect 7681 7759 7691 8041
rect 8123 7759 8133 8041
rect 10911 7663 11343 8041
rect 179 6247 611 6907
rect 3399 6625 3831 7285
rect 3935 6625 4367 7285
rect 7155 7003 7587 7663
rect 7691 7003 8123 7663
rect 10901 7381 10911 7663
rect 11343 7381 11353 7663
rect 10911 6907 11343 7285
rect 179 5491 611 6151
rect 3399 5869 3831 6529
rect 3935 5869 4367 6529
rect 7155 6247 7587 6907
rect 7691 6529 8123 6907
rect 10901 6625 10911 6907
rect 11343 6625 11353 6907
rect 7681 6247 7691 6529
rect 8123 6247 8133 6529
rect 10911 6151 11343 6529
rect 179 4735 611 5395
rect 3399 5113 3831 5773
rect 3935 5113 4367 5773
rect 7155 5491 7587 6151
rect 7691 5773 8123 6151
rect 10901 5869 10911 6151
rect 11343 5869 11353 6151
rect 7681 5491 7691 5773
rect 8123 5491 8133 5773
rect 10911 5395 11343 5773
rect 179 3979 611 4639
rect 3399 4357 3831 5017
rect 3935 4357 4367 5017
rect 7155 4735 7587 5395
rect 7691 5017 8123 5395
rect 10901 5113 10911 5395
rect 11343 5113 11353 5395
rect 7681 4735 7691 5017
rect 8123 4735 8133 5017
rect 10911 4639 11343 5017
rect 3399 3979 4367 4261
rect 7155 3979 7587 4639
rect 7691 4261 8123 4639
rect 10901 4357 10911 4639
rect 11343 4357 11353 4639
rect 7681 3979 7691 4261
rect 8123 3979 8133 4261
rect 10911 3883 11343 4261
rect 179 3223 611 3883
rect 3399 3601 4367 3883
rect 7155 3601 8123 3883
rect 10901 3601 10911 3883
rect 11343 3601 11353 3883
rect 3399 3223 4367 3505
rect 7155 3223 8123 3505
rect 179 2467 611 3127
rect 3399 2845 4367 3127
rect 7155 2845 8123 3127
rect 10911 2845 11343 3505
rect 3399 2467 4367 2749
rect 7155 2467 8123 2749
rect 179 1711 611 2371
rect 3399 2089 4367 2371
rect 7155 2089 8123 2371
rect 10911 2089 11343 2749
rect 3399 1711 4367 1993
rect 7155 1711 8123 1993
rect 179 955 611 1615
rect 3399 1333 4367 1615
rect 7155 1333 8123 1615
rect 10911 1333 11343 1993
rect 3399 955 4367 1237
rect 7155 955 8123 1237
rect 179 199 611 859
rect 3399 577 4367 859
rect 7155 577 8123 859
rect 10911 577 11343 1237
rect 3399 199 4367 481
rect 7155 199 8123 481
rect 10901 199 10911 481
rect 11343 199 11353 481
rect 11447 103 12561 17587
rect -1039 -179 12561 103
rect 12889 477 12961 489
rect 12889 -99 12899 477
rect 12951 -99 12961 477
rect 12889 -111 12961 -99
rect 13011 289 13511 561
rect 13011 89 13161 289
rect 13361 89 13511 289
rect -357 -543 11879 -179
rect 13011 -189 13511 89
rect 13561 6 13789 489
rect 13927 156 13937 222
rect 14003 156 14013 222
rect 13561 -67 14153 6
rect 13561 -111 13860 -67
rect 13585 -543 13860 -111
rect -1259 -791 13860 -543
rect -1259 -1191 -357 -791
rect 14080 -1191 14153 -67
rect -1259 -1438 14153 -1191
<< via1 >>
rect 10921 18253 11333 19108
rect 10911 17209 11343 17491
rect 10911 11161 11343 11443
rect 10911 10405 11343 10687
rect 10911 9649 11343 9931
rect 10911 8893 11343 9175
rect 7691 8515 8123 8797
rect 7691 7759 8123 8041
rect 10911 7381 11343 7663
rect 10911 6625 11343 6907
rect 7691 6247 8123 6529
rect 10911 5869 11343 6151
rect 7691 5491 8123 5773
rect 10911 5113 11343 5395
rect 7691 4735 8123 5017
rect 10911 4357 11343 4639
rect 7691 3979 8123 4261
rect 10911 3601 11343 3883
rect 10911 199 11343 481
rect 12899 -99 12951 477
rect 13161 89 13361 289
rect 13937 131 14003 247
<< metal2 >>
rect 10901 19108 11353 19128
rect 10901 18253 10921 19108
rect 11333 18253 11353 19108
rect 10901 17491 11353 18253
rect 10901 17209 10911 17491
rect 11343 17209 11353 17491
rect 10901 17199 11353 17209
rect 10901 11443 13083 11453
rect 10901 11161 10911 11443
rect 11343 11161 13083 11443
rect 10901 11151 13083 11161
rect 10901 10687 13083 10697
rect 10901 10405 10911 10687
rect 11343 10405 13083 10687
rect 10901 10395 13083 10405
rect 10901 9931 13083 9941
rect 10901 9649 10911 9931
rect 11343 9649 13083 9931
rect 10901 9639 13083 9649
rect 10901 9175 13083 9185
rect 10901 8893 10911 9175
rect 11343 8893 13083 9175
rect 10901 8883 13083 8893
rect 7681 8797 13083 8807
rect 7681 8515 7691 8797
rect 8123 8515 13083 8797
rect 7681 8505 13083 8515
rect 7681 8041 13083 8051
rect 7681 7759 7691 8041
rect 8123 7759 13083 8041
rect 7681 7749 13083 7759
rect 10901 7663 13083 7673
rect 10901 7381 10911 7663
rect 11343 7381 13083 7663
rect 10901 7371 13083 7381
rect 10901 6907 13083 6917
rect 10901 6625 10911 6907
rect 11343 6625 13083 6907
rect 10901 6615 13083 6625
rect 7681 6529 13083 6539
rect 7681 6247 7691 6529
rect 8123 6247 13083 6529
rect 7681 6237 13083 6247
rect 10901 6151 13083 6161
rect 10901 5869 10911 6151
rect 11343 5869 13083 6151
rect 10901 5859 13083 5869
rect 7681 5773 13083 5783
rect 7681 5491 7691 5773
rect 8123 5491 13083 5773
rect 7681 5481 13083 5491
rect 10901 5395 13083 5405
rect 10901 5113 10911 5395
rect 11343 5113 13083 5395
rect 10901 5103 13083 5113
rect 7681 5017 13083 5027
rect 7681 4735 7691 5017
rect 8123 4735 13083 5017
rect 7681 4725 13083 4735
rect 10901 4639 13083 4649
rect 10901 4357 10911 4639
rect 11343 4357 13083 4639
rect 10901 4347 13083 4357
rect 7681 4261 13083 4271
rect 7681 3979 7691 4261
rect 8123 3979 13083 4261
rect 7681 3969 13083 3979
rect 10901 3883 13083 3893
rect 10901 3601 10911 3883
rect 11343 3601 13083 3883
rect 10901 3591 13083 3601
rect 10901 481 12961 491
rect 10901 199 10911 481
rect 11343 477 12961 481
rect 11343 199 12899 477
rect 10901 189 12899 199
rect 12889 -99 12899 189
rect 12951 -99 12961 477
rect 13151 289 14080 299
rect 13151 89 13161 289
rect 13361 247 14080 289
rect 13361 131 13937 247
rect 14003 131 14080 247
rect 13361 89 14080 131
rect 13151 79 14080 89
rect 12889 -111 12961 -99
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 paramcells
timestamp 1713221383
transform 1 0 13970 0 1 189
box -183 -208 183 208
use sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8  sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8_0 paramcells
timestamp 1713221383
transform 1 0 13261 0 1 189
box -528 -558 528 558
use sky130_fd_pr__res_xhigh_po_1p41_H3F4MM  sky130_fd_pr__res_xhigh_po_1p41_H3F4MM_0 paramcells
timestamp 1713221383
transform 0 -1 5761 1 0 8845
box -9024 -5582 9024 5582
use sky130_fd_pr__res_xhigh_po_1p41_LV9PDH  sky130_fd_pr__res_xhigh_po_1p41_LV9PDH_0 paramcells
timestamp 1713221383
transform 0 -1 -482 1 0 8845
box -9024 -557 9024 557
use sky130_fd_pr__res_xhigh_po_1p41_LV9PDH  sky130_fd_pr__res_xhigh_po_1p41_LV9PDH_2
timestamp 1713221383
transform 0 -1 12004 1 0 8845
box -9024 -557 9024 557
<< labels >>
flabel metal1 -1259 18480 -859 18880 3 FreeSans 3200 0 -1200 0 avdd
port 1 e
flabel metal2 12781 3591 13083 3893 3 FreeSans 1280 0 -800 0 out_1111
port 17 e
flabel metal2 12781 3969 13083 4271 3 FreeSans 1280 0 -800 0 out_1110
port 16 e
flabel metal2 12781 4347 13083 4649 3 FreeSans 1280 0 -800 0 out_1101
port 15 e
flabel metal2 12781 4725 13083 5027 3 FreeSans 1280 0 -800 0 out_1100
port 14 e
flabel metal2 12781 5103 13083 5405 3 FreeSans 1280 0 -800 0 out_1011
port 13 e
flabel metal2 12781 5481 13083 5783 3 FreeSans 1280 0 -800 0 out_1010
port 12 e
flabel metal2 12781 5859 13083 6161 3 FreeSans 1280 0 -800 0 out_1001
port 11 e
flabel metal2 12781 6237 13083 6539 3 FreeSans 1280 0 -800 0 out_1000
port 10 e
flabel metal2 12781 6615 13083 6917 3 FreeSans 1280 0 -800 0 out_0111
port 9 e
flabel metal2 12781 7371 13083 7673 3 FreeSans 1280 0 -800 0 out_0110
port 8 e
flabel metal2 12781 7749 13083 8051 3 FreeSans 1280 0 -800 0 out_0101
port 7 e
flabel metal2 12781 8505 13083 8807 3 FreeSans 1280 0 -800 0 out_0100
port 6 e
flabel metal2 12781 8883 13083 9185 3 FreeSans 1280 0 -800 0 out_0011
port 5 e
flabel metal2 12781 9639 13083 9941 3 FreeSans 1280 0 -800 0 out_0010
port 4 e
flabel metal2 12781 10395 13083 10697 3 FreeSans 1280 0 -800 0 out_0001
port 3 e
flabel metal2 12781 11151 13083 11453 3 FreeSans 1280 0 -800 0 out_0000
port 2 e
flabel metal2 13860 79 14080 299 0 FreeSans 1280 0 0 0 ena
port 19 nsew
flabel metal1 7709 11555 8106 11805 0 FreeSans 1280 0 0 0 51
flabel via1 10928 17225 11325 17475 0 FreeSans 1280 0 0 0 138
flabel pwell 7172 17225 7569 17475 0 FreeSans 1280 0 0 0 137
flabel pwell 3416 17225 3813 17475 0 FreeSans 1280 0 0 0 136
flabel pwell 197 16847 594 17097 0 FreeSans 1280 0 0 0 135
flabel pwell 3416 16469 3813 16719 0 FreeSans 1280 0 0 0 134
flabel pwell 197 16091 594 16341 0 FreeSans 1280 0 0 0 133
flabel pwell 3416 15713 3813 15963 0 FreeSans 1280 0 0 0 132
flabel pwell 197 15335 594 15585 0 FreeSans 1280 0 0 0 131
flabel pwell 3416 14957 3813 15207 0 FreeSans 1280 0 0 0 130
flabel pwell 197 14579 594 14829 0 FreeSans 1280 0 0 0 129
flabel pwell 3416 14201 3813 14451 0 FreeSans 1280 0 0 0 128
flabel pwell 197 13823 594 14073 0 FreeSans 1280 0 0 0 127
flabel pwell 3416 13445 3813 13695 0 FreeSans 1280 0 0 0 126
flabel pwell 197 13067 594 13317 0 FreeSans 1280 0 0 0 125
flabel pwell 3416 12689 3813 12939 0 FreeSans 1280 0 0 0 124
flabel pwell 197 12311 594 12561 0 FreeSans 1280 0 0 0 123
flabel pwell 3416 11933 3813 12183 0 FreeSans 1280 0 0 0 122
flabel pwell 197 11555 594 11805 0 FreeSans 1280 0 0 0 121
flabel pwell 3416 11177 3813 11427 0 FreeSans 1280 0 0 0 120
flabel pwell 197 10799 594 11049 0 FreeSans 1280 0 0 0 119
flabel pwell 3416 10421 3813 10671 0 FreeSans 1280 0 0 0 118
flabel pwell 197 10043 594 10293 0 FreeSans 1280 0 0 0 117
flabel pwell 3416 9665 3813 9915 0 FreeSans 1280 0 0 0 116
flabel pwell 197 9287 594 9537 0 FreeSans 1280 0 0 0 115
flabel pwell 3416 8909 3813 9159 0 FreeSans 1280 0 0 0 114
flabel pwell 197 8531 594 8781 0 FreeSans 1280 0 0 0 113
flabel pwell 3416 8153 3813 8403 0 FreeSans 1280 0 0 0 112
flabel pwell 197 7775 594 8025 0 FreeSans 1280 0 0 0 111
flabel pwell 3416 7397 3813 7647 0 FreeSans 1280 0 0 0 110
flabel pwell 197 7019 594 7269 0 FreeSans 1280 0 0 0 109
flabel pwell 3416 6641 3813 6891 0 FreeSans 1280 0 0 0 108
flabel pwell 197 6263 594 6513 0 FreeSans 1280 0 0 0 107
flabel pwell 3416 5885 3813 6135 0 FreeSans 1280 0 0 0 106
flabel pwell 197 5507 594 5757 0 FreeSans 1280 0 0 0 105
flabel pwell 3416 5129 3813 5379 0 FreeSans 1280 0 0 0 104
flabel pwell 197 4751 594 5001 0 FreeSans 1280 0 0 0 103
flabel pwell 3416 4373 3813 4623 0 FreeSans 1280 0 0 0 102
flabel pwell 197 3995 594 4245 0 FreeSans 1280 0 0 0 101
flabel pwell 3953 3995 4350 4245 0 FreeSans 1280 0 0 0 100
flabel pwell 7172 4373 7569 4623 0 FreeSans 1280 0 0 0 99
flabel pwell 3953 4751 4350 5001 0 FreeSans 1280 0 0 0 98
flabel pwell 7172 5129 7569 5379 0 FreeSans 1280 0 0 0 97
flabel pwell 3953 5507 4350 5757 0 FreeSans 1280 0 0 0 96
flabel pwell 7172 5885 7569 6135 0 FreeSans 1280 0 0 0 95
flabel pwell 3953 6263 4350 6513 0 FreeSans 1280 0 0 0 94
flabel pwell 7172 6641 7569 6891 0 FreeSans 1280 0 0 0 93
flabel pwell 3953 7019 4350 7269 0 FreeSans 1280 0 0 0 92
flabel pwell 7172 7397 7569 7647 0 FreeSans 1280 0 0 0 91
flabel pwell 3953 7775 4350 8025 0 FreeSans 1280 0 0 0 90
flabel pwell 7172 8153 7569 8403 0 FreeSans 1280 0 0 0 89
flabel pwell 3953 8531 4350 8781 0 FreeSans 1280 0 0 0 88
flabel pwell 7172 8909 7569 9159 0 FreeSans 1280 0 0 0 87
flabel pwell 3953 9287 4350 9537 0 FreeSans 1280 0 0 0 86
flabel pwell 7172 9665 7569 9915 0 FreeSans 1280 0 0 0 85
flabel pwell 3953 10043 4350 10293 0 FreeSans 1280 0 0 0 84
flabel pwell 7172 10421 7569 10671 0 FreeSans 1280 0 0 0 83
flabel pwell 3953 10799 4350 11049 0 FreeSans 1280 0 0 0 82
flabel pwell 7172 11177 7569 11427 0 FreeSans 1280 0 0 0 81
flabel pwell 3953 11555 4350 11805 0 FreeSans 1280 0 0 0 80
flabel pwell 7172 11933 7569 12183 0 FreeSans 1280 0 0 0 79
flabel pwell 3953 12311 4350 12561 0 FreeSans 1280 0 0 0 78
flabel pwell 7172 12689 7569 12939 0 FreeSans 1280 0 0 0 77
flabel pwell 3953 13067 4350 13317 0 FreeSans 1280 0 0 0 76
flabel pwell 7172 13445 7569 13695 0 FreeSans 1280 0 0 0 75
flabel pwell 3953 13823 4350 14073 0 FreeSans 1280 0 0 0 74
flabel pwell 7172 14201 7569 14451 0 FreeSans 1280 0 0 0 73
flabel pwell 3953 14579 4350 14829 0 FreeSans 1280 0 0 0 72
flabel pwell 7172 14957 7569 15207 0 FreeSans 1280 0 0 0 71
flabel pwell 3953 15335 4350 15585 0 FreeSans 1280 0 0 0 70
flabel pwell 3953 16091 4350 16341 0 FreeSans 1280 0 0 0 68
flabel pwell 7172 15713 7569 15963 0 FreeSans 1280 0 0 0 69
flabel pwell 7172 16469 7569 16719 0 FreeSans 1280 0 0 0 67
flabel pwell 3953 16847 4350 17097 0 FreeSans 1280 0 0 0 66
flabel pwell 10928 16469 11325 16719 0 FreeSans 1280 0 0 0 64
flabel pwell 10928 15713 11325 15963 0 FreeSans 1280 0 0 0 62
flabel pwell 10928 14957 11325 15207 0 FreeSans 1280 0 0 0 60
flabel pwell 10928 14201 11325 14451 0 FreeSans 1280 0 0 0 58
flabel pwell 10928 13445 11325 13695 0 FreeSans 1280 0 0 0 56
flabel pwell 10928 12689 11325 12939 0 FreeSans 1280 0 0 0 54
flabel pwell 10928 11932 11325 12182 0 FreeSans 1280 0 0 0 52
flabel pwell 7709 16847 8106 17097 0 FreeSans 1280 0 0 0 65
flabel pwell 7709 16091 8106 16341 0 FreeSans 1280 0 0 0 63
flabel pwell 7709 15335 8106 15585 0 FreeSans 1280 0 0 0 61
flabel pwell 7709 14579 8106 14829 0 FreeSans 1280 0 0 0 59
flabel pwell 7709 13823 8106 14073 0 FreeSans 1280 0 0 0 57
flabel pwell 7709 13067 8106 13317 0 FreeSans 1280 0 0 0 55
flabel pwell 7709 12311 8106 12561 0 FreeSans 1280 0 0 0 53
flabel pwell 10928 11177 11325 11427 0 FreeSans 1280 0 0 0 50
flabel pwell 7709 10799 8106 11049 0 FreeSans 1280 0 0 0 49
flabel pwell 10928 10421 11325 10671 0 FreeSans 1280 0 0 0 48
flabel pwell 7709 10043 8106 10293 0 FreeSans 1280 0 0 0 47
flabel pwell 10928 9665 11325 9915 0 FreeSans 1280 0 0 0 46
flabel pwell 7709 9287 8106 9537 0 FreeSans 1280 0 0 0 45
flabel pwell 10928 8909 11325 9159 0 FreeSans 1280 0 0 0 44
flabel pwell 7709 8531 8106 8781 0 FreeSans 1280 0 0 0 43
flabel pwell 10928 8153 11325 8403 0 FreeSans 1280 0 0 0 42
flabel pwell 7709 7775 8106 8025 0 FreeSans 1280 0 0 0 41
flabel pwell 10928 7397 11325 7647 0 FreeSans 1280 0 0 0 40
flabel pwell 7709 7019 8106 7269 0 FreeSans 1280 0 0 0 39
flabel pwell 10928 6641 11325 6891 0 FreeSans 1280 0 0 0 38
flabel pwell 7709 6263 8106 6513 0 FreeSans 1280 0 0 0 37
flabel pwell 10928 5885 11325 6135 0 FreeSans 1280 0 0 0 36
flabel pwell 7709 5507 8106 5757 0 FreeSans 1280 0 0 0 35
flabel pwell 10928 5129 11325 5379 0 FreeSans 1280 0 0 0 34
flabel pwell 7709 4751 8106 5001 0 FreeSans 1280 0 0 0 33
flabel pwell 10928 4373 11325 4623 0 FreeSans 1280 0 0 0 32
flabel pwell 7709 3995 8106 4245 0 FreeSans 1280 0 0 0 31
flabel pwell 10928 3617 11325 3867 0 FreeSans 1280 0 0 0 30
flabel pwell 7172 3617 7569 3867 0 FreeSans 1280 0 0 0 29
flabel pwell 3416 3617 3813 3867 0 FreeSans 1280 0 0 0 28
flabel pwell 197 3239 594 3489 0 FreeSans 1280 0 0 0 27
flabel pwell 3953 3239 4350 3489 0 FreeSans 1280 0 0 0 26
flabel pwell 7709 3239 8106 3489 0 FreeSans 1280 0 0 0 25
flabel pwell 10928 2861 11325 3111 0 FreeSans 1280 0 0 0 24
flabel pwell 7172 2861 7569 3111 0 FreeSans 1280 0 0 0 23
flabel pwell 3416 2861 3813 3111 0 FreeSans 1280 0 0 0 22
flabel pwell 197 2483 594 2733 0 FreeSans 1280 0 0 0 21
flabel pwell 3953 2483 4350 2733 0 FreeSans 1280 0 0 0 20
flabel pwell 7709 2483 8106 2733 0 FreeSans 1280 0 0 0 19
flabel pwell 10928 2105 11325 2355 0 FreeSans 1280 0 0 0 18
flabel pwell 7172 2105 7569 2355 0 FreeSans 1280 0 0 0 17
flabel pwell 3416 2105 3813 2355 0 FreeSans 1280 0 0 0 16
flabel pwell 197 1727 594 1977 0 FreeSans 1280 0 0 0 15
flabel pwell 3953 1727 4350 1977 0 FreeSans 1280 0 0 0 14
flabel pwell 7709 1727 8106 1977 0 FreeSans 1280 0 0 0 13
flabel pwell 10928 1349 11325 1599 0 FreeSans 1280 0 0 0 12
flabel pwell 7172 1349 7569 1599 0 FreeSans 1280 0 0 0 11
flabel pwell 3416 1349 3813 1599 0 FreeSans 1280 0 0 0 10
flabel pwell 197 971 594 1221 0 FreeSans 1280 0 0 0 9
flabel pwell 3953 971 4350 1221 0 FreeSans 1280 0 0 0 8
flabel pwell 7709 971 8106 1221 0 FreeSans 1280 0 0 0 7
flabel pwell 10928 593 11325 843 0 FreeSans 1280 0 0 0 6
flabel pwell 7172 593 7569 843 0 FreeSans 1280 0 0 0 5
flabel pwell 3416 593 3813 843 0 FreeSans 1280 0 0 0 4
flabel pwell 197 215 594 465 0 FreeSans 1280 0 0 0 3
flabel pwell 3953 215 4350 465 0 FreeSans 1280 0 0 0 2
flabel pwell 7709 215 8106 465 0 FreeSans 1280 0 0 0 1
flabel metal1 -1259 -1191 -859 -791 3 FreeSans 3200 0 -1200 0 avss
port 18 e
<< properties >>
string MASKHINTS_HVI -1248 17909 12770 18077 -1248 -388 12770 -220
<< end >>
